// From https://github.com/icebreaker-fpga/icebreaker-workshop
// Seven segment controller
// Switches quickly between the two parts of the display
// to create the illusion of both halves being illuminated
// at the same time.
module seven_seg_ctrl (
    input CLK,
    input [7:0] din,
    output reg [7:0] dout
);
    wire [6:0] lsb_digit;
    wire [6:0] msb_digit;

    seven_seg_hex msb_nibble (
        .din(din[7:4]),
        .dout(msb_digit)
    );

    seven_seg_hex lsb_nibble (
        .din(din[3:0]),
        .dout(lsb_digit)
    );

    reg [9:0] clkdiv = 0;
    reg clkdiv_pulse = 0;
    reg msb_not_lsb = 0;

    always @(posedge CLK) begin
        clkdiv <= clkdiv + 1;
        clkdiv_pulse <= &clkdiv;
        msb_not_lsb <= msb_not_lsb ^ clkdiv_pulse;

        if (clkdiv_pulse) begin
            if (msb_not_lsb) begin
                dout[6:0] <= ~msb_digit;
                dout[7] <= 0;
            end else begin
                dout[6:0] <= ~lsb_digit;
                dout[7] <= 1;
            end
        end
    end
endmodule

// From https://github.com/icebreaker-fpga/icebreaker-workshop
// Convert 4bit numbers to 7 segments
module seven_seg_hex (
    input [3:0] din,
    output reg [6:0] dout
);
    always @*
        case (din)
            4'h0: dout = 7'b 0111111;
            4'h1: dout = 7'b 0000110;
            4'h2: dout = 7'b 1011011;
            4'h3: dout = 7'b 1001111;
            4'h4: dout = 7'b 1100110;
            4'h5: dout = 7'b 1101101;
            4'h6: dout = 7'b 1111101;
            4'h7: dout = 7'b 0000111;
            4'h8: dout = 7'b 1111111;
            4'h9: dout = 7'b 1101111;
            4'hA: dout = 7'b 1110111;
            4'hB: dout = 7'b 1111100;
            4'hC: dout = 7'b 0111001;
            4'hD: dout = 7'b 1011110;
            4'hE: dout = 7'b 1111001;
            4'hF: dout = 7'b 1110001;
            default: dout = 7'b 1000000;
        endcase
endmodule